module ROB(
    port_list
);
  
endmodule