`timescale 1ps/1ps;
`include "../common/micro_op.svh"


module free_list_tb;
  


endmodule