//////////////////////////////////////////////////////////////////////////////////
// Project Name: RIA
// Create Date: 2021/06/08
// Contributor: Jian Shi
// Reviewer: 
// Module Name: rob
// Target Devices: reorder buffer
// Description: 
// track the state of all inflight instructions in the pipeline
// Dependencies: 
// src/common/micro_op.svh, src/frontend/rat.sv
//////////////////////////////////////////////////////////////////////////////////
`include "../common/micro_op.svh"

module rob (
  input     clock
);
  
endmodule
