// Project: RISC-V SoC Microarchitecture Design & Optimization
// Module:  Ria (Top Module)
// Author:  Li Shi
// Date:    2021/06/21

