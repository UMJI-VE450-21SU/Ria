`ifndef __DEFINES_SVH__
`define __DEFINES_SVH__



`endif  // __DEFINES_SVH__
